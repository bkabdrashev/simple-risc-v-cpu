localparam RS =  473630 ;
